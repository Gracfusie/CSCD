// -----------------------------------------------------------------------------
// Memory-like top wrapper for the PE core.
// - 32-bit word port matches the simple SRAM-like slave used in the lab setup.
// - No wait states; reads return registered data in 1 cycle.
// Map this block to a base address (e.g., 0x7000_0000) via the AXI crossbar,
// and bridge with axi2mem like SRAM (see lab example).  :contentReference[oaicite:3]{index=3}
// -----------------------------------------------------------------------------
module NPU_top #(
  parameter int N = 10,
  parameter int K_SIZE = 3,
  parameter int DATA_WIDTH = 8,
  parameter int AXI_WIDTH = 32,
  parameter int ADDR_W = 3  // enough for 0..4
) (
  input  logic               clk,
  input  logic               rst_n,        // high-active

  // SRAM-like memory port (compatible with axi2mem style)
  input  logic               req_i,        // access qualifier (assume always 1'b1 OK)
  input  logic [3:0]         wen_i,        // byte enables; write if any bit=1
  input  logic [ADDR_W-1:0]  addr_i,       // word index (offset / 4)
  input  logic [AXI_WIDTH-1:0]        wdata_i,
  output logic [AXI_WIDTH-1:0]        rdata_o
);

  // NPU buffer
  parameter int BUFFER_DEPTH = (2*N+1)*K_SIZE;          // 63
  parameter int SEL_DEMUX_WIDTH = $clog2(BUFFER_DEPTH); // 6
  logic [K_SIZE*DATA_WIDTH-1:0] npu_buffer [0:BUFFER_DEPTH-1];
  logic [DATA_WIDTH-1:0] npu_buffer_flattened [0:K_SIZE*BUFFER_DEPTH-1];
  always_comb begin
    for (int i = 0; i < BUFFER_DEPTH; i++) begin
      for (int j = 0; j < K_SIZE; j++) begin
        npu_buffer_flattened[i*K_SIZE + j] = npu_buffer[i][(j+1)*DATA_WIDTH-1 -: DATA_WIDTH];
      end
    end
  end
  // assign npu_buffer_flattened = npu_buffer;

  // MUX parameters
  parameter int MUX_A_DEPTH = K_SIZE*K_SIZE;           // 9
  parameter int SEL_MUX_A_WIDTH = $clog2(MUX_A_DEPTH); // 4
  parameter int MUX_B_DEPTH = K_SIZE*K_SIZE*2;         // 18
  parameter int SEL_MUX_B_WIDTH = $clog2(MUX_B_DEPTH); // 5

  // NPU scheduler
  wire [N-1:0] pe_en, pe_mode_sel, pe_reg_reset;
  wire [SEL_DEMUX_WIDTH-1:0] pe_demux_sel;
  wire [SEL_MUX_A_WIDTH-1:0] pe_mux_a_sel;
  wire [SEL_MUX_B_WIDTH-1:0] pe_mux_b_sel;
  npu_scheduler #(
    .N               (N),
    .W_IN            (DATA_WIDTH),
    .SEL_DEMUX_WIDTH (SEL_DEMUX_WIDTH),
    .SEL_MUX_A_WIDTH (SEL_MUX_A_WIDTH),
    .SEL_MUX_B_WIDTH (SEL_MUX_B_WIDTH)
  ) u_npu_scheduler (
    .clk          (clk),
    .rst_n        (rst_n),
    .instr        (wdata_i[AXI_WIDTH-1:AXI_WIDTH-DATA_WIDTH]),

    .pe_en        (pe_en),
    .pe_mode_sel  (pe_mode_sel),
    .pe_reg_reset (pe_reg_reset),
    .pe_demux_sel (pe_demux_sel),
    .pe_mux_a_sel (pe_mux_a_sel),
    .pe_mux_b_sel (pe_mux_b_sel)
  );

  // Write demux
  // (0-9)*9 for weights, (10-19)*9 for direct inputs, 20*9 for broadcast inputs
  wire [BUFFER_DEPTH*K*DATA_WIDTH-1:0] npu_buffer_wdata;
  wire [BUFFER_DEPTH-1:0] npu_buffer_wen;

  pe_demux #(
    .DATA_WIDTH (K_SIZE*DATA_WIDTH),
    .DATA_DEPTH (BUFFER_DEPTH),
    .SEL_WIDTH  (SEL_DEMUX_WIDTH)
  ) u_demux (
    .data_in (wdata_i[K_SIZE*DATA_WIDTH-1:0]),
    .sel     (pe_demux_sel),
    .en      (|wen_i),
    .data_out(npu_buffer_wdata)
  );

  pe_binary_decoder #(
    .ADDR_WIDTH (SEL_DEMUX_WIDTH),
    .DEPTH      (BUFFER_DEPTH)
  ) u_decoder (
    .addr (pe_demux_sel),
    .en   (|wen_i),
    .y    (npu_buffer_wen)
  );

  always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      for (int i = 0; i < BUFFER_DEPTH; i++) begin
        npu_buffer[i] <= '0;
      end
      rdata_o <= '0;
    end else begin
      // Write operation
      for (int i = 0; i < BUFFER_DEPTH; i++) begin
        if (npu_buffer_wen[i]) begin
          npu_buffer[i] <= npu_buffer_wdata[(i+1)*(K_SIZE*DATA_WIDTH)-1 -: K_SIZE*DATA_WIDTH];
        end
      end
    end    
  end

  // Read mux
  wire [DATA_WIDTH-1:0] a_mul [N-1:0];
  wire [DATA_WIDTH-1:0] b_mul [N-1:0];

  generate
    for (genvar i = 0; i < N; i++) begin : PE_MUX_GEN_WEIGHT
      pe_mux #(
        .WIDTH     (DATA_WIDTH),
        .DEPTH     (MUX_A_DEPTH),
        .SEL_WIDTH (SEL_MUX_A_WIDTH)
      ) u_pe_mux (
        .data_in (npu_buffer_flattened[i*MUX_A_DEPTH +: MUX_A_DEPTH]),
        .sel     (pe_mux_a_sel),
        .data_out(a_mul[i])
      );
    end
  endgenerate

  generate
    for (genvar i = 0; i < N; i++) begin : PE_MUX_GEN_INPUT
      wire [DATA_WIDTH-1:0] data_in [0:MUX_B_DEPTH-1];
      assign data_in[0:MUX_A_DEPTH-1] = npu_buffer_flattened[(N+i)*MUX_A_DEPTH +: MUX_A_DEPTH];
      assign data_in[MUX_A_DEPTH:MUX_B_DEPTH-1] = npu_buffer_flattened[2*N*MUX_A_DEPTH +: MUX_A_DEPTH];

      pe_mux #(
        .WIDTH    (DATA_WIDTH),
        .DEPTH    (MUX_B_DEPTH),
        .SEL_WIDTH(SEL_MUX_B_WIDTH)
      ) u_pe_mux (
        // .data_in ({npu_buffer_flattened[(N+i)*MUX_A_DEPTH +: MUX_A_DEPTH], npu_buffer_flattened[2*N*MUX_A_DEPTH +: MUX_A_DEPTH]}),
        .data_in (data_in),
        .sel     (pe_mux_b_sel),
        .data_out(b_mul[i])
      );
    end
  endgenerate

  // PE cores
  generate
    for (genvar i = 0; i < N; i++) begin: PE_CORE_GEN
      pe_core #(
        .W_IN (DATA_WIDTH),
        .W_MUL(2*DATA_WIDTH),
        .W_ACC(3*DATA_WIDTH)
      ) u_pe_core (
        .clk      (clk),
        .rst_n    (rst_n),
        .pe_en    (pe_en[i]),
        .mode_sel (pe_mode_sel[i]),
        .reg_reset(pe_reg_reset[i]),
        .a_mul     (a_mul[i]),
        .b_mul     (b_mul[i]),
        .results  ()
      );
    end
  endgenerate



endmodule
